module main;
	initial begin
		$display("Hello World!\n");
	end
endmodule
module half_adder(input wire a, input wire b, output wire sum, output wire carry);
	assign sum = a^b;
	assign carry = a&b;
endmodule

// https://i.sstatic.net/E0itr.png
module full_adder(input wire a, input wire b, input wire in_carry, output wire sum, output wire out_carry);
	wire first_add;
	wire [1:0] half_adder_carries;

	half_adder ha0 ( 
		.a(a),
		.b(b),
		.sum(first_add),
		.carry(half_adder_carries[0])
	);
	half_adder ha1 (
		.a(first_add),
		.b(in_carry),
		.sum(sum),
		.carry(half_adder_carries[1])
	);
	assign out_carry = half_adder_carries[0]|half_adder_carries[1];
endmodule

module adder #(parameter WIDTH = 8) (
	input wire [WIDTH-1:0] a,
	input wire [WIDTH-1:0] b,
	output wire [WIDTH-1:0] sum,
	output wire overflow
);
	wire [WIDTH-1:0] adder_carries;
	half_adder ha (
		.a(a[0]),
		.b(b[0]),
		.sum(sum[0]),
		.carry(adder_carries[0])
	);

	genvar i;
	generate
		for(i = 1; i < WIDTH; i = i + 1) begin: adder_loop
			full_adder fa (
				.a(a[i]),
				.b(b[i]),
				.in_carry(adder_carries[i-1]),
				.sum(sum[i]),
				.out_carry(adder_carries[i])
			);
		end
	endgenerate

	assign overflow = adder_carries[WIDTH-1];
endmodule

module main;
 	reg [3:0] a;
	reg [3:0] b;
	wire [3:0] sum;
	wire overflow; 

 
	adder #(.WIDTH(4)) uut (
		.a(a),
		.b(b),
		.sum(sum),
		.overflow(overflow)
	);

	initial begin
        $monitor("[Time: %0d]\t%b + %b = %b\t(overflow=%b)\n", $time, a, b, sum, overflow);
		a = 4'b0111; b = 4'b1101; #10; // 7 - 3 = 4 (sign bit on left)
		a = 4'b1001; b = 4'b1111; #10; // -7 - 1 = -8 
        $finish;    
	end
endmodule